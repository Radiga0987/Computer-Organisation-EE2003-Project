//Module for all control signals of the accelerator
module control_mm(       
	input opcode_1
	input 


);